[{"type":"Conceptual","source_relative_path":"articles/glossary.md","output":{".html":{"relative_path":"articles/glossary.html","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX\\obj\\.cache\\build\\ufdwnla1.opp\\dzoaqeg1.urj","hash":"zf+ghQp7g6Os2OUH0NgoJoFcMjwq4SCMhdpLSEvkWpc="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"glossary\" sourcefile=\"articles/glossary.md\" sourcestartlinenumber=\"1\">Glossary</h1>"},{"type":"Conceptual","source_relative_path":"articles/application-hierarchy.md","output":{".html":{"relative_path":"articles/application-hierarchy.html","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX\\obj\\.cache\\build\\ufdwnla1.opp\\x051iyo3.qfd","hash":"xMm7fKL354ODfdLKyw0nrBef8Rk5+yBSnxTPy+X4Htg="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"application-hierarchy-and-interitence\" sourcefile=\"articles/application-hierarchy.md\" sourcestartlinenumber=\"1\">Application Hierarchy and Interitence</h1>"},{"type":"Conceptual","source_relative_path":"articles/create-application-using-hyperconsole.md","output":{".html":{"relative_path":"articles/create-application-using-hyperconsole.html","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX\\obj\\.cache\\build\\ufdwnla1.opp\\t32p4ecp.kfz","hash":"KPqfdH/Xl0NcDRgHhAgfJ4Jtp2LDYKRUHe1e5xEs2Ms="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"create-application-using-hyperconsole\" sourcefile=\"articles/create-application-using-hyperconsole.md\" sourcestartlinenumber=\"1\">Create Application Using Hyperconsole</h1>"},{"type":"Conceptual","source_relative_path":"README.md","output":{".html":{"relative_path":"README.html","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX\\obj\\.cache\\build\\ufdwnla1.opp\\dg31rmd1.km2","hash":"/4qGEroixst7Ed902o30zw/ZjkdhMMje1ODdo0c3gXU="}},"is_incremental":true,"version":"","rawTitle":"<h2 id=\"description\" sourcefile=\"README.md\" sourcestartlinenumber=\"1\">Description</h2>"},{"type":"Conceptual","source_relative_path":"api/index.md","output":{".html":{"relative_path":"api/index.html","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX\\obj\\.cache\\build\\ufdwnla1.opp\\vaqrhrkn.0zo","hash":"wszsSMPYzapVndH8Qeyv7cB01DhHFSiHKSiE4OBzeh8="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"placeholder\" sourcefile=\"api/index.md\" sourcestartlinenumber=\"1\">PLACEHOLDER</h1>"},{"type":"Conceptual","source_relative_path":"articles/create-application-introduction.md","output":{".html":{"relative_path":"articles/create-application-introduction.html","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX\\obj\\.cache\\build\\ufdwnla1.opp\\atbyxqoc.xzw","hash":"qaLM2lnK9+4flWAh0szgwyyvezOgIabHIfYFYnC/9sI="}},"is_incremental":false,"version":"","rawTitle":"<h1 id=\"create-application\" sourcefile=\"articles/create-application-introduction.md\" sourcestartlinenumber=\"1\">Create Application</h1>"},{"type":"Toc","source_relative_path":"api/toc.yml","output":{".html":{"relative_path":"api/toc.html","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX\\obj\\.cache\\build\\ufdwnla1.opp\\kcxgldig.m0l","hash":"53cDPdjyKTmYSaPMwcMYYJO/bYpeY21eGi/JWyVQBqE="}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.8New.png","output":{"resource":{"relative_path":"articles/resources/2.8New.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.8New.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.16DeleteAppSearch.png","output":{"resource":{"relative_path":"articles/resources/2.16DeleteAppSearch.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.16DeleteAppSearch.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/emgage-logo-large-transparent-2.png","output":{"resource":{"relative_path":"articles/resources/emgage-logo-large-transparent-2.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/emgage-logo-large-transparent-2.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/4.Search.png","output":{"resource":{"relative_path":"articles/resources/4.Search.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/4.Search.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.11-PublishDraftApp.png","output":{"resource":{"relative_path":"articles/resources/2.11-PublishDraftApp.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.11-PublishDraftApp.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.10-FindAndPublish.png","output":{"resource":{"relative_path":"articles/resources/2.10-FindAndPublish.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.10-FindAndPublish.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/Screenshot 2022-09-22 190721.png","output":{"resource":{"relative_path":"articles/resources/Screenshot 2022-09-22 190721.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/Screenshot 2022-09-22 190721.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.9-Launch.png","output":{"resource":{"relative_path":"articles/resources/2.9-Launch.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.9-Launch.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.14DiscardDraft.png","output":{"resource":{"relative_path":"articles/resources/2.14DiscardDraft.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.14DiscardDraft.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/1.1login.png","output":{"resource":{"relative_path":"articles/resources/1.1login.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/1.1login.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/images/logo.png","output":{"resource":{"relative_path":"articles/images/logo.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/images/logo.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.7New.png","output":{"resource":{"relative_path":"articles/resources/2.7New.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.7New.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.1Dashboard-Search.png","output":{"resource":{"relative_path":"articles/resources/2.1Dashboard-Search.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.1Dashboard-Search.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/1.2login.png","output":{"resource":{"relative_path":"articles/resources/1.2login.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/1.2login.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.19PUblishInside.png","output":{"resource":{"relative_path":"articles/resources/2.19PUblishInside.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.19PUblishInside.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.13PublishDraft.png","output":{"resource":{"relative_path":"articles/resources/2.13PublishDraft.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.13PublishDraft.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.16DEleteAppClear.png","output":{"resource":{"relative_path":"articles/resources/2.16DEleteAppClear.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.16DEleteAppClear.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.15DiscardDraftInside.png","output":{"resource":{"relative_path":"articles/resources/2.15DiscardDraftInside.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.15DiscardDraftInside.png"}},"is_incremental":false,"version":""},{"type":"Toc","source_relative_path":"articles/toc.yml","output":{".html":{"relative_path":"articles/toc.html","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX\\obj\\.cache\\build\\ufdwnla1.opp\\nzyqupvj.jmi","hash":"AJzhOjJmRJdjG9axE6amHak/9ZcLo9syn9kXUMYpMM8="}},"is_incremental":false,"version":""},{"type":"Toc","source_relative_path":"toc.yml","output":{".html":{"relative_path":"toc.html","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX\\obj\\.cache\\build\\ufdwnla1.opp\\ztazcrij.gpa","hash":"vNoj18SCkAxmWuMVrvurDfDS+LocAZOZiirN4I0GYiw="}},"is_incremental":false,"version":""},{"type":"Conceptual","source_relative_path":"articles/create-application-using-appmanager.md","output":{".html":{"relative_path":"articles/create-application-using-appmanager.html","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX\\obj\\.cache\\build\\ufdwnla1.opp\\qfv5evl2.g05","hash":"PT9XPQ7AJTEn060wbchoMNydKMSPOw3BKaJeczbRc44="}},"is_incremental":false,"version":"","rawTitle":"<h1 id=\"create-application-using-app-manager\" sourcefile=\"articles/create-application-using-appmanager.md\" sourcestartlinenumber=\"1\">Create Application Using App Manager</h1>"},{"type":"Conceptual","source_relative_path":"articles/articles-introduction.md","output":{".html":{"relative_path":"articles/articles-introduction.html","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX\\obj\\.cache\\build\\ufdwnla1.opp\\34njpmp3.4a0","hash":"MwZ3vM/eBqZY2VPgBoM8U6GiL5FD34X/rP0NhcYMGFk="}},"is_incremental":false,"version":"","rawTitle":"<h1 id=\"emgage-documentation\" sourcefile=\"articles/articles-introduction.md\" sourcestartlinenumber=\"1\">Emgage Documentation</h1>"},{"type":"Resource","source_relative_path":"articles/resources/1.png","output":{"resource":{"relative_path":"articles/resources/1.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/1.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.1New.png","output":{"resource":{"relative_path":"articles/resources/2.1New.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.1New.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/1.4login.png","output":{"resource":{"relative_path":"articles/resources/1.4login.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/1.4login.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.6New.png","output":{"resource":{"relative_path":"articles/resources/2.6New.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.6New.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.5New.png","output":{"resource":{"relative_path":"articles/resources/2.5New.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.5New.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.2New-Publish.png","output":{"resource":{"relative_path":"articles/resources/2.2New-Publish.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.2New-Publish.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/1.login.png","output":{"resource":{"relative_path":"articles/resources/1.login.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/1.login.png"}},"is_incremental":false,"version":""},{"type":"Conceptual","source_relative_path":"index.md","output":{".html":{"relative_path":"index.html","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX\\obj\\.cache\\build\\ufdwnla1.opp\\gkdqxofe.2fo","hash":"Yahic1gvH5Id1OGbSyUjxt6RtlcqksLitrodsiaWNOA="}},"is_incremental":false,"version":"","rawTitle":"<h2 id=\"about-emgage\" sourcefile=\"index.md\" sourcestartlinenumber=\"1\">About Emgage</h2>"},{"type":"Resource","source_relative_path":"articles/resources/Screenshot 2022-09-22 190428.png","output":{"resource":{"relative_path":"articles/resources/Screenshot 2022-09-22 190428.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/Screenshot 2022-09-22 190428.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/emgage-squarelogo-1469225763276.png","output":{"resource":{"relative_path":"articles/resources/emgage-squarelogo-1469225763276.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/emgage-squarelogo-1469225763276.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.19DeleteInside.png","output":{"resource":{"relative_path":"articles/resources/2.19DeleteInside.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.19DeleteInside.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.3New.png","output":{"resource":{"relative_path":"articles/resources/2.3New.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.3New.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.2New.png","output":{"resource":{"relative_path":"articles/resources/2.2New.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.2New.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/3.3Editsettings.png","output":{"resource":{"relative_path":"articles/resources/3.3Editsettings.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/3.3Editsettings.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.Dashboard.png","output":{"resource":{"relative_path":"articles/resources/2.Dashboard.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.Dashboard.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.12-DeleteAnApp.png","output":{"resource":{"relative_path":"articles/resources/2.12-DeleteAnApp.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.12-DeleteAnApp.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/3.Hyperconsole-New.png","output":{"resource":{"relative_path":"articles/resources/3.Hyperconsole-New.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/3.Hyperconsole-New.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.1Dashboard-Clear.png","output":{"resource":{"relative_path":"articles/resources/2.1Dashboard-Clear.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.1Dashboard-Clear.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/4.Search-clear.png","output":{"resource":{"relative_path":"articles/resources/4.Search-clear.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/4.Search-clear.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.12-DeleteAnApp - Copy.png","output":{"resource":{"relative_path":"articles/resources/2.12-DeleteAnApp - Copy.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.12-DeleteAnApp - Copy.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"articles/resources/2.13PublishDraftClear.png","output":{"resource":{"relative_path":"articles/resources/2.13PublishDraftClear.png","link_to_path":"D:\\zHammadHassan\\UpWork\\001.Emgage\\02-Contract02\\EmgageDocFX/articles/resources/2.13PublishDraftClear.png"}},"is_incremental":false,"version":""}]